yvyyyggyyy