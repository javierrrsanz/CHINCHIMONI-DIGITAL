ijfidfijfjefeifdefijndfjednf
hola buenas tardes
