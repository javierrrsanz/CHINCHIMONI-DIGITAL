ijfidfijfjefeifdefijndfjednf